library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

-- A 128x8 single-port RAM in VHDL
entity memory is
port(
 RAM_ADDR: in std_logic_vector(15 downto 0); -- Address to write/read RAM
 RAM_DATA_IN: in std_logic_vector(15 downto 0); -- Data to write into RAM
 RAM_WR: in std_logic; -- Write enable 
 RAM_CLOCK: in std_logic; -- clock input for RAM
 RAM_DATA_OUT: out std_logic_vector(15 downto 0) -- Data output of RAM
);
end memory;

architecture Behavioral of memory is
-- define the new type for the 65535x16 RAM 
type RAM_ARRAY is array (0 to  65535) of std_logic_vector (15 downto 0);
-- initial values in the RAM
signal RAM: RAM_ARRAY :=(
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
	   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"5555",x"6666",x"7777",x"6767",-- 0x00: 
   x"9999",x"0000",x"0000",x"1111",-- 0x04: 
   x"0000",x"0000",x"0000",x"0000",-- 0x08: 
   x"0000",x"0000",x"0000",x"0000",-- 0x0C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x10: 
   x"0000",x"0000",x"0000",x"0000",-- 0x14: 
   x"0000",x"0000",x"0000",x"0000",-- 0x18: 
   x"0000",x"0000",x"0000",x"0000",-- 0x1C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x20: 
   x"0000",x"0000",x"0000",x"0000",-- 0x24: 
   x"0000",x"0000",x"0000",x"0000",-- 0x28: 
   x"0000",x"0000",x"0000",x"0000",-- 0x2C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x30: 
   x"0000",x"0000",x"0000",x"0000",-- 0x34: 
   x"0000",x"0000",x"0000",x"0000",-- 0x38: 
   x"0000",x"0000",x"0000",x"0000",-- 0x3C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x40: 
   x"0000",x"0000",x"0000",x"0000",-- 0x44: 
   x"0000",x"0000",x"0000",x"0000",-- 0x48: 
   x"0000",x"0000",x"0000",x"0000",-- 0x4C: 
   x"0000",x"0000",x"0000",x"0000",-- 0x50: 
   x"0000",x"0000",x"0000",x"0000",-- 0x54: 
   x"0000",x"0000",x"0000",x"0000",-- 0x58: 
   x"0000",x"0000",x"0000",x"0000",-- 0x5C: 
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000",
   x"0000",x"0000",x"0000",x"0000"

   ); 
begin
process(RAM_CLOCK)
begin
 if(rising_edge(RAM_CLOCK)) then
 if(RAM_WR='1') then -- when write enable = 1, 
 -- write input data into RAM at the provided address
 RAM(to_integer(unsigned(RAM_ADDR))) <= RAM_DATA_IN;
 -- The index of the RAM array type needs to be integer so
 -- converts RAM_ADDR from std_logic_vector -> Unsigned -> Interger using numeric_std library
 end if;
 end if;
end process;
 -- Data to be read out 
 RAM_DATA_OUT <= RAM(to_integer(unsigned(RAM_ADDR)));
end Behavioral;
